/*
Problem statement: Implement the following circuit:
                    output always ground 
                    
Solution:
*/

module top_module (
    output out);
assign out= 1'b0;
endmodule
