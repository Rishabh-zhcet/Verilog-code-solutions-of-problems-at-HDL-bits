/*
Problem Statement: Implement the following circuit:
                    in--------> out
                    
Solution:

*/

module top_module (
    input in,
    output out);
    
    assign out=in;

endmodule

