// Problem statement: Build a circuit with no inputs and one output. That output should always drive 1 (or logic high).

//Solution:

module top_module( output wire one );

    assign one =1;

endmodule
